module test #(input logic param = 4)(
    input foo,
    input bar
);

function automatic foo();
  return;
endfunction

logic [2:0] a = "foo";
logic bar[4] = foo;
logic another[bar] = foo;
logic another bar[r]
logic another bar[3:0];

  LOCALPARAM a = 3;

endmodule
